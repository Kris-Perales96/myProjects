module ALU_tb;

reg aluOF, aluCarry, enable, clk, reset;
reg[7:0] aluSum, A, B;
reg [3:0] opcode;

PowerALU_Kristopher_Perales alu1(aluSum,, aluCarry, aluOF, enable, opcode, A, B, clk, reset);

initial
begin
	reset = 1'b1;
	clk = 1'b0;
	forever #10 clk = ~clk;
	forever #30 reset = ~reset;
end

initial
begin
	opcode = 4'd0;
	forever #10 opcode = opcode + 1;
end

initial
begin
   #20 A = 8'b10011001; B = 4'b1001000;
   #20 A = 8'b10011000; B = 4'b1001010;
   #20 A = 8'b10011101; B = 4'b1001111;
   #20 A = 8'b10010100; B = 4'b1001100;
   #20 A = 8'b10010101; B = 4'b1001010;
   #20 A = 8'b10010001; B = 4'b1001100;
   #20 A = 8'b10011111; B = 4'b1001101;
   #20 A = 8'b10011010; B = 4'b1001000;
   #20 A = 8'b10010111; B = 4'b1001111;
   #20 A = 8'b10011010; B = 4'b1001110;
   #20 A = 8'b10011000; B = 4'b1001011;
   #20 A = 8'b10011010; B = 4'b1001111;
   #20 A = 8'b10011000; B = 4'b1001011;
   #20 A = 8'b10011011; B = 4'b1001101;
   #20 A = 8'b10011000; B = 4'b1001100;
   #20 A = 8'b10011111; B = 4'b1001010;
   #20 A = 8'b10010011; B = 4'b1001111;
   #20 A = 8'b10010001; B = 4'b1001001;
   #20 A = 8'b10010001; B = 4'b1001001;
   #20 A = 8'b10010001; B = 4'b1001000;
   #20 A = 8'b10010110; B = 4'b1001101;
   #20 A = 8'b10010111; B = 4'b1001100;
   #20 A = 8'b10010101; B = 4'b1001110;
   #20 A = 8'b10011100; B = 4'b1001011;
   #20 A = 8'b10011010; B = 4'b1001111;
   #20 A = 8'b10011100; B = 4'b1001110;
   #20 A = 8'b10011110; B = 4'b1001100;
   #20 A = 8'b10011111; B = 4'b1001000;
   #20 A = 8'b10010011; B = 4'b1001010;
   #20 A = 8'b10010010; B = 4'b1001100;
   #20 A = 8'b10011011; B = 4'b1001011;
   #20 A = 8'b10010001; B = 4'b1001000;
   #20 A = 8'b10011000; B = 4'b1001100;
   #20 A = 8'b10011000; B = 4'b1001100;
   #20 A = 8'b10011101; B = 4'b1001011;
   #20 A = 8'b10010111; B = 4'b1001001;
   #20 A = 8'b10010110; B = 4'b1001111;
   #20 A = 8'b10011010; B = 4'b1001110;
   #20 A = 8'b10011011; B = 4'b1001100;
   #20 A = 8'b10011000; B = 4'b1001010;
   #20 A = 8'b10010101; B = 4'b1001000;
   #20 A = 8'b10010010; B = 4'b1001010;
   #20 A = 8'b10011001; B = 4'b1001000;
   #20 A = 8'b10010100; B = 4'b1001001;
   #20 A = 8'b10010000; B = 4'b1001010;
   #20 A = 8'b10011100; B = 4'b1001000;
   #20 A = 8'b10010011; B = 4'b1001010;
   #20 A = 8'b10010111; B = 4'b1001000;
   #20 A = 8'b10011011; B = 4'b1001001;
   #20 A = 8'b10010101; B = 4'b1001111;
   #20 A = 8'b10011011; B = 4'b1001100;
   #20 A = 8'b10010110; B = 4'b1001000;
   #20 A = 8'b10011010; B = 4'b1001111;
   #20 A = 8'b10011011; B = 4'b1001011;
   #20 A = 8'b10010111; B = 4'b1001011;
   #20 A = 8'b10010000; B = 4'b1001000;
   #20 A = 8'b10010101; B = 4'b1001111;
   #20 A = 8'b10010110; B = 4'b1001101;
   #20 A = 8'b10010100; B = 4'b1001011;
   #20 A = 8'b10010011; B = 4'b1001011;
   #20 A = 8'b10011101; B = 4'b1001001;
   #20 A = 8'b10010110; B = 4'b1001000;
   #20 A = 8'b10011110; B = 4'b1001000;
   #20 A = 8'b10010110; B = 4'b1001010;
   #20 A = 8'b10011100; B = 4'b1001110;
   #20 A = 8'b10010110; B = 4'b1001101;
   #20 A = 8'b10011100; B = 4'b1001111;
   #20 A = 8'b10011100; B = 4'b1001000;
   #20 A = 8'b10010110; B = 4'b1001101;
   #20 A = 8'b10010011; B = 4'b1001000;
   #20 A = 8'b10011100; B = 4'b1001001;
   #20 A = 8'b10011111; B = 4'b1001000;
   #20 A = 8'b10010101; B = 4'b1001101;
   #20 A = 8'b10011010; B = 4'b1001101;
   #20 A = 8'b10010111; B = 4'b1001000;
   #20 A = 8'b10011101; B = 4'b1001010;
   #20 A = 8'b10011100; B = 4'b1001101;
   #20 A = 8'b10010010; B = 4'b1001101;
   #20 A = 8'b10011101; B = 4'b1001110;
   #20 A = 8'b10011111; B = 4'b1001010;
   #20 A = 8'b10011000; B = 4'b1001111;
   #20 A = 8'b10011110; B = 4'b1001010;
   #20 A = 8'b10011001; B = 4'b1001100;
   #20 A = 8'b10010010; B = 4'b1001101;
   #20 A = 8'b10010011; B = 4'b1001010;
   #20 A = 8'b10010110; B = 4'b1001010;
   #20 A = 8'b10011011; B = 4'b1001110;
   #20 A = 8'b10011101; B = 4'b1001001;
   #20 A = 8'b10011100; B = 4'b1001011;
   #20 A = 8'b10010101; B = 4'b1001100;
   #20 A = 8'b10011000; B = 4'b1001111;
   #20 A = 8'b10010001; B = 4'b1001000;
   #20 A = 8'b10010001; B = 4'b1001101;
end

endmodule
